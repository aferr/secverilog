module quant_ternary_vqe();
//-----------------------------------------------------------------------------
// Ternary operators
//-----------------------------------------------------------------------------
wire [3:0] {L} a;
wire [3:0] {|i| Par 1 ? 0 : 1} b;

//sat
assign a[0] = b[0];
//unsat
assign a[0] = b[1];

endmodule
