module arrtype();

reg[1:0] { |i| a | b} foo;


endmodule
