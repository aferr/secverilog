module quant_boolean();
wire [3:0] {L} a;
wire [3:0] {|i| Par (3==4)} b;

endmodule
