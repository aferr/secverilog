module quant_basic();


   //-----------------------------------------------------------------------------
   // Ignore non-index
   //-----------------------------------------------------------------------------
   wire [1:0] {L} a;

   wire [1:0] {|i| LH 0} b;


   //should pass
   assign a[0] = b[0];

   //should pass
   assign a[1] = b[1];


   //-----------------------------------------------------------------------------
   // Use index
   //-----------------------------------------------------------------------------
   wire [1:0] {L} c;

   wire [1:0] {|i| LH i} d;


   //should pass
   assign c[0] = d[0];

   //should fail
   assign c[1] = d[1];


   //-----------------------------------------------------------------------------
   // Quantifying over indexing expression (1)
   //-----------------------------------------------------------------------------
   wire [1:0] {L} e;

   wire [1:0] {|i| LH i} f;

   wire       g;


   //should fail
   assign e[0] = f[g];


   //-----------------------------------------------------------------------------
   // Quantifying over indexing expression (2)
   //-----------------------------------------------------------------------------
   wire [1:0] {L} h;

   wire [1:0] {|i| LH 0} i;

   wire       j;


   //should pass
   assign h[0] = i[j];


   //-----------------------------------------------------------------------------
   // Quantifying over indexing expression (3)
   //-----------------------------------------------------------------------------
   wire [1:0] {|i| LH i} k;

   wire [1:0] {|i| LH i} l;


   //should pass
   assign k[0] = l[0];

   //should pass
   assign k[1] = l[1];


   //-----------------------------------------------------------------------------
   // Quantified Join Types (1)
   //-----------------------------------------------------------------------------
   wire [1:0] {|i| LH i} m;

   wire [1:0] {|i| LH i} n;

   wire [1:0] {H} o;


   //should fail
   assign m[0] = n[0] + o[0];

   //should pass
   assign m[1] = n[1] + o[1];


   //-----------------------------------------------------------------------------
   // Quantified Join Types (1)
   //-----------------------------------------------------------------------------
   wire [1:0] {|i| LH i} p;

   wire [1:0] {|i| LH i} q;

   wire [1:0] {|i| LH i} r;


   //should pass
   assign p[0] = q[0] + r[0];

   //should pass
   assign p[1] = q[1] + r[1];


endmodule
